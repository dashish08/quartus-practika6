library verilog;
use verilog.vl_types.all;
entity practika6_vlg_vec_tst is
end practika6_vlg_vec_tst;
